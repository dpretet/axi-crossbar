`ifndef TB_FUNCTIONS
`define TB_FUNCTIONS
function automatic integer gen_resp(integer data);

    gen_resp = ~data;

endfunction
`endif
